library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ram_contrasenas is
	port(data0,data1,data2,data3,data4: in std_logic_vector(3 downto 0);
	add: in std_logic_vector(3 downto 0);
	modo,reset: in std_logic;
	t0,t1,t2,t3,t4: buffer std_logic_vector(3 downto 0);--fija
	q0,q1,q2,q3,q4: buffer std_logic_vector(3 downto 0));--variable
end ram_contrasenas;
architecture sol of ram_contrasenas is
signal r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,cualquiera: std_logic_vector(3 downto 0);
signal r10,r11,r12,r13,r14,r15,r16,r17,r18,r19: std_logic_vector(3 downto 0);
signal r20,r21,r22,r23,r24,r25,r26,r27,r28,r29: std_logic_vector(3 downto 0);
signal r30,r31,r32,r33,r34,r35,r36,r37,r38,r39: std_logic_vector(3 downto 0);
signal r40,r41,r42,r43,r44,r45,r46,r47,r48,r49: std_logic_vector(3 downto 0);
begin
		process(modo,add)
			begin
				if reset='0' then r45<="0000";t0<="0000";
						r46<="0001";t1<="0001";
						r47<="0010";t2<="0010";
						r48<="0011";t3<="0011";
						r49<="0100";t4<="0100";
				elsif modo='1' then --escritura
					case add is
						when "0000" => r0<=data0;
						r1<=data1;
						r2<=data2;
						r3<=data3;
						r4<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "0001" =>r5<=data0;
						r6<=data1;
						r7<=data2;
						r8<=data3;
						r9<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "0010" => r10<=data0;
						r11<=data1;
						r12<=data2;
						r13<=data3;
						r14<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "0011" => r15<=data0;
						r16<=data1;
						r17<=data2;
						r18<=data3;
						r19<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "0100" => r20<=data0;
						r21<=data1;
						r22<=data2;
						r23<=data3;
						r24<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "0101" => r25<=data0;
						r26<=data1;
						r27<=data2;
						r28<=data3;
						r29<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "0110" => r30<=data0;
						r31<=data1;
						r32<=data2;
						r33<=data3;
						r34<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "0111" => r35<=data0;
						r36<=data1;
						r37<=data2;
						r38<=data3;
						r39<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "1000" => r40<=data0;
						r41<=data1;
						r42<=data2;
						r43<=data3;
						r44<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when "1001" => r45<=data0;
						r46<=data1;
						r47<=data2;
						r48<=data3;
						r49<=data4;
						t0<=data0;
						t1<=data1;
						t2<=data2;
						t3<=data3;
						t4<=data4;
						when others => cualquiera<="0000";
					end case;
				
				else
					case add is--lectura
						when "0000" => q0<=r0;
						q1<=r1;
						q2<=r2;
						q3<=r3;
						q4<=r4;
						when "0001" => q0<=r5;
						q1<=r6;
						q2<=r7;
						q3<=r8;
						q4<=r9;
						when "0010" => q0<=r10;
						q1<=r11;
						q2<=r12;
						q3<=r13;
						q4<=r14;
						when "0011" => q0<=r15;
						q1<=r16;
						q2<=r17;
						q3<=r18;
						q4<=r19;
						when "0100" => q0<=r20;
						q1<=r21;
						q2<=r22;
						q3<=r23;
						q4<=r24;
						when "0101" => q0<=r25;
						q1<=r26;
						q2<=r27;
						q3<=r28;
						q4<=r29;
						when "0110" => q0<=r30;
						q1<=r31;
						q2<=r32;
						q3<=r33;
						q4<=r34;
						when "0111" => q0<=r35;
						q1<=r36;
						q2<=r37;
						q3<=r38;
						q4<=r39;
						when "1000" => q0<=r40;
						q1<=r41;
						q2<=r42;
						q3<=r43;
						q4<=r44;
						when "1001" => q0<=r45;
						q1<=r46;
						q2<=r47;
						q3<=r48;
						q4<=r49;
						when others => cualquiera<="0000";
					end case;
				end if;
	end process;
end sol;